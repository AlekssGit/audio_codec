library verilog;
use verilog.vl_types.all;
entity audio_codec is
    port(
        clock           : in     vl_logic
    );
end audio_codec;
